// For 512-point IFFT
// 8 read ports

module ifft_twiddle_rom (
  input [7:0] addr0,
  input [7:0] addr1,
  input [7:0] addr2,
  input [7:0] addr3,
  input [7:0] addr4,
  input [7:0] addr5,
  input [7:0] addr6,
  input [7:0] addr7,
  output [15:0] data0_re,
  output [15:0] data0_im,
  output [15:0] data1_re,
  output [15:0] data1_im,
  output [15:0] data2_re,
  output [15:0] data2_im,
  output [15:0] data3_re,
  output [15:0] data3_im,
  output [15:0] data4_re,
  output [15:0] data4_im,
  output [15:0] data5_re,
  output [15:0] data5_im,
  output [15:0] data6_re,
  output [15:0] data6_im,
  output [15:0] data7_re,
  output [15:0] data7_im
);
  // For N=512
  wire signed [15:0] wn_re [0:255];
  wire signed [15:0] wn_im [0:255];

  assign wn_re[0] = $signed(16'sh7FFF);
  assign wn_re[1] = $signed(16'sh7FFE);
  assign wn_re[2] = $signed(16'sh7FF6);
  assign wn_re[3] = $signed(16'sh7FEA);
  assign wn_re[4] = $signed(16'sh7FD9);
  assign wn_re[5] = $signed(16'sh7FC2);
  assign wn_re[6] = $signed(16'sh7FA7);
  assign wn_re[7] = $signed(16'sh7F87);
  assign wn_re[8] = $signed(16'sh7F62);
  assign wn_re[9] = $signed(16'sh7F38);
  assign wn_re[10] = $signed(16'sh7F0A);
  assign wn_re[11] = $signed(16'sh7ED6);
  assign wn_re[12] = $signed(16'sh7E9D);
  assign wn_re[13] = $signed(16'sh7E60);
  assign wn_re[14] = $signed(16'sh7E1E);
  assign wn_re[15] = $signed(16'sh7DD6);
  assign wn_re[16] = $signed(16'sh7D8A);
  assign wn_re[17] = $signed(16'sh7D3A);
  assign wn_re[18] = $signed(16'sh7CE4);
  assign wn_re[19] = $signed(16'sh7C89);
  assign wn_re[20] = $signed(16'sh7C2A);
  assign wn_re[21] = $signed(16'sh7BC6);
  assign wn_re[22] = $signed(16'sh7B5D);
  assign wn_re[23] = $signed(16'sh7AEF);
  assign wn_re[24] = $signed(16'sh7A7D);
  assign wn_re[25] = $signed(16'sh7A06);
  assign wn_re[26] = $signed(16'sh798A);
  assign wn_re[27] = $signed(16'sh790A);
  assign wn_re[28] = $signed(16'sh7885);
  assign wn_re[29] = $signed(16'sh77FB);
  assign wn_re[30] = $signed(16'sh776C);
  assign wn_re[31] = $signed(16'sh76D9);
  assign wn_re[32] = $signed(16'sh7642);
  assign wn_re[33] = $signed(16'sh75A6);
  assign wn_re[34] = $signed(16'sh7505);
  assign wn_re[35] = $signed(16'sh7460);
  assign wn_re[36] = $signed(16'sh73B6);
  assign wn_re[37] = $signed(16'sh7308);
  assign wn_re[38] = $signed(16'sh7255);
  assign wn_re[39] = $signed(16'sh719E);
  assign wn_re[40] = $signed(16'sh70E3);
  assign wn_re[41] = $signed(16'sh7023);
  assign wn_re[42] = $signed(16'sh6F5F);
  assign wn_re[43] = $signed(16'sh6E97);
  assign wn_re[44] = $signed(16'sh6DCA);
  assign wn_re[45] = $signed(16'sh6CF9);
  assign wn_re[46] = $signed(16'sh6C24);
  assign wn_re[47] = $signed(16'sh6B4B);
  assign wn_re[48] = $signed(16'sh6A6E);
  assign wn_re[49] = $signed(16'sh698C);
  assign wn_re[50] = $signed(16'sh68A7);
  assign wn_re[51] = $signed(16'sh67BD);
  assign wn_re[52] = $signed(16'sh66D0);
  assign wn_re[53] = $signed(16'sh65DE);
  assign wn_re[54] = $signed(16'sh64E9);
  assign wn_re[55] = $signed(16'sh63EF);
  assign wn_re[56] = $signed(16'sh62F2);
  assign wn_re[57] = $signed(16'sh61F1);
  assign wn_re[58] = $signed(16'sh60EC);
  assign wn_re[59] = $signed(16'sh5FE4);
  assign wn_re[60] = $signed(16'sh5ED7);
  assign wn_re[61] = $signed(16'sh5DC8);
  assign wn_re[62] = $signed(16'sh5CB4);
  assign wn_re[63] = $signed(16'sh5B9D);
  assign wn_re[64] = $signed(16'sh5A82);
  assign wn_re[65] = $signed(16'sh5964);
  assign wn_re[66] = $signed(16'sh5843);
  assign wn_re[67] = $signed(16'sh571E);
  assign wn_re[68] = $signed(16'sh55F6);
  assign wn_re[69] = $signed(16'sh54CA);
  assign wn_re[70] = $signed(16'sh539B);
  assign wn_re[71] = $signed(16'sh5269);
  assign wn_re[72] = $signed(16'sh5134);
  assign wn_re[73] = $signed(16'sh4FFB);
  assign wn_re[74] = $signed(16'sh4EC0);
  assign wn_re[75] = $signed(16'sh4D81);
  assign wn_re[76] = $signed(16'sh4C40);
  assign wn_re[77] = $signed(16'sh4AFB);
  assign wn_re[78] = $signed(16'sh49B4);
  assign wn_re[79] = $signed(16'sh486A);
  assign wn_re[80] = $signed(16'sh471D);
  assign wn_re[81] = $signed(16'sh45CD);
  assign wn_re[82] = $signed(16'sh447B);
  assign wn_re[83] = $signed(16'sh4326);
  assign wn_re[84] = $signed(16'sh41CE);
  assign wn_re[85] = $signed(16'sh4074);
  assign wn_re[86] = $signed(16'sh3F17);
  assign wn_re[87] = $signed(16'sh3DB8);
  assign wn_re[88] = $signed(16'sh3C57);
  assign wn_re[89] = $signed(16'sh3AF3);
  assign wn_re[90] = $signed(16'sh398D);
  assign wn_re[91] = $signed(16'sh3825);
  assign wn_re[92] = $signed(16'sh36BA);
  assign wn_re[93] = $signed(16'sh354E);
  assign wn_re[94] = $signed(16'sh33DF);
  assign wn_re[95] = $signed(16'sh326E);
  assign wn_re[96] = $signed(16'sh30FC);
  assign wn_re[97] = $signed(16'sh2F87);
  assign wn_re[98] = $signed(16'sh2E11);
  assign wn_re[99] = $signed(16'sh2C99);
  assign wn_re[100] = $signed(16'sh2B1F);
  assign wn_re[101] = $signed(16'sh29A4);
  assign wn_re[102] = $signed(16'sh2827);
  assign wn_re[103] = $signed(16'sh26A8);
  assign wn_re[104] = $signed(16'sh2528);
  assign wn_re[105] = $signed(16'sh23A7);
  assign wn_re[106] = $signed(16'sh2224);
  assign wn_re[107] = $signed(16'sh209F);
  assign wn_re[108] = $signed(16'sh1F1A);
  assign wn_re[109] = $signed(16'sh1D93);
  assign wn_re[110] = $signed(16'sh1C0C);
  assign wn_re[111] = $signed(16'sh1A83);
  assign wn_re[112] = $signed(16'sh18F9);
  assign wn_re[113] = $signed(16'sh176E);
  assign wn_re[114] = $signed(16'sh15E2);
  assign wn_re[115] = $signed(16'sh1455);
  assign wn_re[116] = $signed(16'sh12C8);
  assign wn_re[117] = $signed(16'sh113A);
  assign wn_re[118] = $signed(16'sh0FAB);
  assign wn_re[119] = $signed(16'sh0E1C);
  assign wn_re[120] = $signed(16'sh0C8C);
  assign wn_re[121] = $signed(16'sh0AFB);
  assign wn_re[122] = $signed(16'sh096B);
  assign wn_re[123] = $signed(16'sh07D9);
  assign wn_re[124] = $signed(16'sh0648);
  assign wn_re[125] = $signed(16'sh04B6);
  assign wn_re[126] = $signed(16'sh0324);
  assign wn_re[127] = $signed(16'sh0192);
  assign wn_re[128] = $signed(16'sh0000);
  assign wn_re[129] = $signed(-16'sh0192);
  assign wn_re[130] = $signed(-16'sh0324);
  assign wn_re[131] = $signed(-16'sh04B6);
  assign wn_re[132] = $signed(-16'sh0648);
  assign wn_re[133] = $signed(-16'sh07D9);
  assign wn_re[134] = $signed(-16'sh096B);
  assign wn_re[135] = $signed(-16'sh0AFB);
  assign wn_re[136] = $signed(-16'sh0C8C);
  assign wn_re[137] = $signed(-16'sh0E1C);
  assign wn_re[138] = $signed(-16'sh0FAB);
  assign wn_re[139] = $signed(-16'sh113A);
  assign wn_re[140] = $signed(-16'sh12C8);
  assign wn_re[141] = $signed(-16'sh1455);
  assign wn_re[142] = $signed(-16'sh15E2);
  assign wn_re[143] = $signed(-16'sh176E);
  assign wn_re[144] = $signed(-16'sh18F9);
  assign wn_re[145] = $signed(-16'sh1A83);
  assign wn_re[146] = $signed(-16'sh1C0C);
  assign wn_re[147] = $signed(-16'sh1D93);
  assign wn_re[148] = $signed(-16'sh1F1A);
  assign wn_re[149] = $signed(-16'sh209F);
  assign wn_re[150] = $signed(-16'sh2224);
  assign wn_re[151] = $signed(-16'sh23A7);
  assign wn_re[152] = $signed(-16'sh2528);
  assign wn_re[153] = $signed(-16'sh26A8);
  assign wn_re[154] = $signed(-16'sh2827);
  assign wn_re[155] = $signed(-16'sh29A4);
  assign wn_re[156] = $signed(-16'sh2B1F);
  assign wn_re[157] = $signed(-16'sh2C99);
  assign wn_re[158] = $signed(-16'sh2E11);
  assign wn_re[159] = $signed(-16'sh2F87);
  assign wn_re[160] = $signed(-16'sh30FC);
  assign wn_re[161] = $signed(-16'sh326E);
  assign wn_re[162] = $signed(-16'sh33DF);
  assign wn_re[163] = $signed(-16'sh354E);
  assign wn_re[164] = $signed(-16'sh36BA);
  assign wn_re[165] = $signed(-16'sh3825);
  assign wn_re[166] = $signed(-16'sh398D);
  assign wn_re[167] = $signed(-16'sh3AF3);
  assign wn_re[168] = $signed(-16'sh3C57);
  assign wn_re[169] = $signed(-16'sh3DB8);
  assign wn_re[170] = $signed(-16'sh3F17);
  assign wn_re[171] = $signed(-16'sh4074);
  assign wn_re[172] = $signed(-16'sh41CE);
  assign wn_re[173] = $signed(-16'sh4326);
  assign wn_re[174] = $signed(-16'sh447B);
  assign wn_re[175] = $signed(-16'sh45CD);
  assign wn_re[176] = $signed(-16'sh471D);
  assign wn_re[177] = $signed(-16'sh486A);
  assign wn_re[178] = $signed(-16'sh49B4);
  assign wn_re[179] = $signed(-16'sh4AFB);
  assign wn_re[180] = $signed(-16'sh4C40);
  assign wn_re[181] = $signed(-16'sh4D81);
  assign wn_re[182] = $signed(-16'sh4EC0);
  assign wn_re[183] = $signed(-16'sh4FFB);
  assign wn_re[184] = $signed(-16'sh5134);
  assign wn_re[185] = $signed(-16'sh5269);
  assign wn_re[186] = $signed(-16'sh539B);
  assign wn_re[187] = $signed(-16'sh54CA);
  assign wn_re[188] = $signed(-16'sh55F6);
  assign wn_re[189] = $signed(-16'sh571E);
  assign wn_re[190] = $signed(-16'sh5843);
  assign wn_re[191] = $signed(-16'sh5964);
  assign wn_re[192] = $signed(-16'sh5A82);
  assign wn_re[193] = $signed(-16'sh5B9D);
  assign wn_re[194] = $signed(-16'sh5CB4);
  assign wn_re[195] = $signed(-16'sh5DC8);
  assign wn_re[196] = $signed(-16'sh5ED7);
  assign wn_re[197] = $signed(-16'sh5FE4);
  assign wn_re[198] = $signed(-16'sh60EC);
  assign wn_re[199] = $signed(-16'sh61F1);
  assign wn_re[200] = $signed(-16'sh62F2);
  assign wn_re[201] = $signed(-16'sh63EF);
  assign wn_re[202] = $signed(-16'sh64E9);
  assign wn_re[203] = $signed(-16'sh65DE);
  assign wn_re[204] = $signed(-16'sh66D0);
  assign wn_re[205] = $signed(-16'sh67BD);
  assign wn_re[206] = $signed(-16'sh68A7);
  assign wn_re[207] = $signed(-16'sh698C);
  assign wn_re[208] = $signed(-16'sh6A6E);
  assign wn_re[209] = $signed(-16'sh6B4B);
  assign wn_re[210] = $signed(-16'sh6C24);
  assign wn_re[211] = $signed(-16'sh6CF9);
  assign wn_re[212] = $signed(-16'sh6DCA);
  assign wn_re[213] = $signed(-16'sh6E97);
  assign wn_re[214] = $signed(-16'sh6F5F);
  assign wn_re[215] = $signed(-16'sh7023);
  assign wn_re[216] = $signed(-16'sh70E3);
  assign wn_re[217] = $signed(-16'sh719E);
  assign wn_re[218] = $signed(-16'sh7255);
  assign wn_re[219] = $signed(-16'sh7308);
  assign wn_re[220] = $signed(-16'sh73B6);
  assign wn_re[221] = $signed(-16'sh7460);
  assign wn_re[222] = $signed(-16'sh7505);
  assign wn_re[223] = $signed(-16'sh75A6);
  assign wn_re[224] = $signed(-16'sh7642);
  assign wn_re[225] = $signed(-16'sh76D9);
  assign wn_re[226] = $signed(-16'sh776C);
  assign wn_re[227] = $signed(-16'sh77FB);
  assign wn_re[228] = $signed(-16'sh7885);
  assign wn_re[229] = $signed(-16'sh790A);
  assign wn_re[230] = $signed(-16'sh798A);
  assign wn_re[231] = $signed(-16'sh7A06);
  assign wn_re[232] = $signed(-16'sh7A7D);
  assign wn_re[233] = $signed(-16'sh7AEF);
  assign wn_re[234] = $signed(-16'sh7B5D);
  assign wn_re[235] = $signed(-16'sh7BC6);
  assign wn_re[236] = $signed(-16'sh7C2A);
  assign wn_re[237] = $signed(-16'sh7C89);
  assign wn_re[238] = $signed(-16'sh7CE4);
  assign wn_re[239] = $signed(-16'sh7D3A);
  assign wn_re[240] = $signed(-16'sh7D8A);
  assign wn_re[241] = $signed(-16'sh7DD6);
  assign wn_re[242] = $signed(-16'sh7E1E);
  assign wn_re[243] = $signed(-16'sh7E60);
  assign wn_re[244] = $signed(-16'sh7E9D);
  assign wn_re[245] = $signed(-16'sh7ED6);
  assign wn_re[246] = $signed(-16'sh7F0A);
  assign wn_re[247] = $signed(-16'sh7F38);
  assign wn_re[248] = $signed(-16'sh7F62);
  assign wn_re[249] = $signed(-16'sh7F87);
  assign wn_re[250] = $signed(-16'sh7FA7);
  assign wn_re[251] = $signed(-16'sh7FC2);
  assign wn_re[252] = $signed(-16'sh7FD9);
  assign wn_re[253] = $signed(-16'sh7FEA);
  assign wn_re[254] = $signed(-16'sh7FF6);
  assign wn_re[255] = $signed(-16'sh7FFE);
  assign wn_im[0] = $signed(16'sh0000);
  assign wn_im[1] = $signed(16'sh0192);
  assign wn_im[2] = $signed(16'sh0324);
  assign wn_im[3] = $signed(16'sh04B6);
  assign wn_im[4] = $signed(16'sh0648);
  assign wn_im[5] = $signed(16'sh07D9);
  assign wn_im[6] = $signed(16'sh096B);
  assign wn_im[7] = $signed(16'sh0AFB);
  assign wn_im[8] = $signed(16'sh0C8C);
  assign wn_im[9] = $signed(16'sh0E1C);
  assign wn_im[10] = $signed(16'sh0FAB);
  assign wn_im[11] = $signed(16'sh113A);
  assign wn_im[12] = $signed(16'sh12C8);
  assign wn_im[13] = $signed(16'sh1455);
  assign wn_im[14] = $signed(16'sh15E2);
  assign wn_im[15] = $signed(16'sh176E);
  assign wn_im[16] = $signed(16'sh18F9);
  assign wn_im[17] = $signed(16'sh1A83);
  assign wn_im[18] = $signed(16'sh1C0C);
  assign wn_im[19] = $signed(16'sh1D93);
  assign wn_im[20] = $signed(16'sh1F1A);
  assign wn_im[21] = $signed(16'sh209F);
  assign wn_im[22] = $signed(16'sh2224);
  assign wn_im[23] = $signed(16'sh23A7);
  assign wn_im[24] = $signed(16'sh2528);
  assign wn_im[25] = $signed(16'sh26A8);
  assign wn_im[26] = $signed(16'sh2827);
  assign wn_im[27] = $signed(16'sh29A4);
  assign wn_im[28] = $signed(16'sh2B1F);
  assign wn_im[29] = $signed(16'sh2C99);
  assign wn_im[30] = $signed(16'sh2E11);
  assign wn_im[31] = $signed(16'sh2F87);
  assign wn_im[32] = $signed(16'sh30FC);
  assign wn_im[33] = $signed(16'sh326E);
  assign wn_im[34] = $signed(16'sh33DF);
  assign wn_im[35] = $signed(16'sh354E);
  assign wn_im[36] = $signed(16'sh36BA);
  assign wn_im[37] = $signed(16'sh3825);
  assign wn_im[38] = $signed(16'sh398D);
  assign wn_im[39] = $signed(16'sh3AF3);
  assign wn_im[40] = $signed(16'sh3C57);
  assign wn_im[41] = $signed(16'sh3DB8);
  assign wn_im[42] = $signed(16'sh3F17);
  assign wn_im[43] = $signed(16'sh4074);
  assign wn_im[44] = $signed(16'sh41CE);
  assign wn_im[45] = $signed(16'sh4326);
  assign wn_im[46] = $signed(16'sh447B);
  assign wn_im[47] = $signed(16'sh45CD);
  assign wn_im[48] = $signed(16'sh471D);
  assign wn_im[49] = $signed(16'sh486A);
  assign wn_im[50] = $signed(16'sh49B4);
  assign wn_im[51] = $signed(16'sh4AFB);
  assign wn_im[52] = $signed(16'sh4C40);
  assign wn_im[53] = $signed(16'sh4D81);
  assign wn_im[54] = $signed(16'sh4EC0);
  assign wn_im[55] = $signed(16'sh4FFB);
  assign wn_im[56] = $signed(16'sh5134);
  assign wn_im[57] = $signed(16'sh5269);
  assign wn_im[58] = $signed(16'sh539B);
  assign wn_im[59] = $signed(16'sh54CA);
  assign wn_im[60] = $signed(16'sh55F6);
  assign wn_im[61] = $signed(16'sh571E);
  assign wn_im[62] = $signed(16'sh5843);
  assign wn_im[63] = $signed(16'sh5964);
  assign wn_im[64] = $signed(16'sh5A82);
  assign wn_im[65] = $signed(16'sh5B9D);
  assign wn_im[66] = $signed(16'sh5CB4);
  assign wn_im[67] = $signed(16'sh5DC8);
  assign wn_im[68] = $signed(16'sh5ED7);
  assign wn_im[69] = $signed(16'sh5FE4);
  assign wn_im[70] = $signed(16'sh60EC);
  assign wn_im[71] = $signed(16'sh61F1);
  assign wn_im[72] = $signed(16'sh62F2);
  assign wn_im[73] = $signed(16'sh63EF);
  assign wn_im[74] = $signed(16'sh64E9);
  assign wn_im[75] = $signed(16'sh65DE);
  assign wn_im[76] = $signed(16'sh66D0);
  assign wn_im[77] = $signed(16'sh67BD);
  assign wn_im[78] = $signed(16'sh68A7);
  assign wn_im[79] = $signed(16'sh698C);
  assign wn_im[80] = $signed(16'sh6A6E);
  assign wn_im[81] = $signed(16'sh6B4B);
  assign wn_im[82] = $signed(16'sh6C24);
  assign wn_im[83] = $signed(16'sh6CF9);
  assign wn_im[84] = $signed(16'sh6DCA);
  assign wn_im[85] = $signed(16'sh6E97);
  assign wn_im[86] = $signed(16'sh6F5F);
  assign wn_im[87] = $signed(16'sh7023);
  assign wn_im[88] = $signed(16'sh70E3);
  assign wn_im[89] = $signed(16'sh719E);
  assign wn_im[90] = $signed(16'sh7255);
  assign wn_im[91] = $signed(16'sh7308);
  assign wn_im[92] = $signed(16'sh73B6);
  assign wn_im[93] = $signed(16'sh7460);
  assign wn_im[94] = $signed(16'sh7505);
  assign wn_im[95] = $signed(16'sh75A6);
  assign wn_im[96] = $signed(16'sh7642);
  assign wn_im[97] = $signed(16'sh76D9);
  assign wn_im[98] = $signed(16'sh776C);
  assign wn_im[99] = $signed(16'sh77FB);
  assign wn_im[100] = $signed(16'sh7885);
  assign wn_im[101] = $signed(16'sh790A);
  assign wn_im[102] = $signed(16'sh798A);
  assign wn_im[103] = $signed(16'sh7A06);
  assign wn_im[104] = $signed(16'sh7A7D);
  assign wn_im[105] = $signed(16'sh7AEF);
  assign wn_im[106] = $signed(16'sh7B5D);
  assign wn_im[107] = $signed(16'sh7BC6);
  assign wn_im[108] = $signed(16'sh7C2A);
  assign wn_im[109] = $signed(16'sh7C89);
  assign wn_im[110] = $signed(16'sh7CE4);
  assign wn_im[111] = $signed(16'sh7D3A);
  assign wn_im[112] = $signed(16'sh7D8A);
  assign wn_im[113] = $signed(16'sh7DD6);
  assign wn_im[114] = $signed(16'sh7E1E);
  assign wn_im[115] = $signed(16'sh7E60);
  assign wn_im[116] = $signed(16'sh7E9D);
  assign wn_im[117] = $signed(16'sh7ED6);
  assign wn_im[118] = $signed(16'sh7F0A);
  assign wn_im[119] = $signed(16'sh7F38);
  assign wn_im[120] = $signed(16'sh7F62);
  assign wn_im[121] = $signed(16'sh7F87);
  assign wn_im[122] = $signed(16'sh7FA7);
  assign wn_im[123] = $signed(16'sh7FC2);
  assign wn_im[124] = $signed(16'sh7FD9);
  assign wn_im[125] = $signed(16'sh7FEA);
  assign wn_im[126] = $signed(16'sh7FF6);
  assign wn_im[127] = $signed(16'sh7FFE);
  assign wn_im[128] = $signed(16'sh7FFF);
  assign wn_im[129] = $signed(16'sh7FFE);
  assign wn_im[130] = $signed(16'sh7FF6);
  assign wn_im[131] = $signed(16'sh7FEA);
  assign wn_im[132] = $signed(16'sh7FD9);
  assign wn_im[133] = $signed(16'sh7FC2);
  assign wn_im[134] = $signed(16'sh7FA7);
  assign wn_im[135] = $signed(16'sh7F87);
  assign wn_im[136] = $signed(16'sh7F62);
  assign wn_im[137] = $signed(16'sh7F38);
  assign wn_im[138] = $signed(16'sh7F0A);
  assign wn_im[139] = $signed(16'sh7ED6);
  assign wn_im[140] = $signed(16'sh7E9D);
  assign wn_im[141] = $signed(16'sh7E60);
  assign wn_im[142] = $signed(16'sh7E1E);
  assign wn_im[143] = $signed(16'sh7DD6);
  assign wn_im[144] = $signed(16'sh7D8A);
  assign wn_im[145] = $signed(16'sh7D3A);
  assign wn_im[146] = $signed(16'sh7CE4);
  assign wn_im[147] = $signed(16'sh7C89);
  assign wn_im[148] = $signed(16'sh7C2A);
  assign wn_im[149] = $signed(16'sh7BC6);
  assign wn_im[150] = $signed(16'sh7B5D);
  assign wn_im[151] = $signed(16'sh7AEF);
  assign wn_im[152] = $signed(16'sh7A7D);
  assign wn_im[153] = $signed(16'sh7A06);
  assign wn_im[154] = $signed(16'sh798A);
  assign wn_im[155] = $signed(16'sh790A);
  assign wn_im[156] = $signed(16'sh7885);
  assign wn_im[157] = $signed(16'sh77FB);
  assign wn_im[158] = $signed(16'sh776C);
  assign wn_im[159] = $signed(16'sh76D9);
  assign wn_im[160] = $signed(16'sh7642);
  assign wn_im[161] = $signed(16'sh75A6);
  assign wn_im[162] = $signed(16'sh7505);
  assign wn_im[163] = $signed(16'sh7460);
  assign wn_im[164] = $signed(16'sh73B6);
  assign wn_im[165] = $signed(16'sh7308);
  assign wn_im[166] = $signed(16'sh7255);
  assign wn_im[167] = $signed(16'sh719E);
  assign wn_im[168] = $signed(16'sh70E3);
  assign wn_im[169] = $signed(16'sh7023);
  assign wn_im[170] = $signed(16'sh6F5F);
  assign wn_im[171] = $signed(16'sh6E97);
  assign wn_im[172] = $signed(16'sh6DCA);
  assign wn_im[173] = $signed(16'sh6CF9);
  assign wn_im[174] = $signed(16'sh6C24);
  assign wn_im[175] = $signed(16'sh6B4B);
  assign wn_im[176] = $signed(16'sh6A6E);
  assign wn_im[177] = $signed(16'sh698C);
  assign wn_im[178] = $signed(16'sh68A7);
  assign wn_im[179] = $signed(16'sh67BD);
  assign wn_im[180] = $signed(16'sh66D0);
  assign wn_im[181] = $signed(16'sh65DE);
  assign wn_im[182] = $signed(16'sh64E9);
  assign wn_im[183] = $signed(16'sh63EF);
  assign wn_im[184] = $signed(16'sh62F2);
  assign wn_im[185] = $signed(16'sh61F1);
  assign wn_im[186] = $signed(16'sh60EC);
  assign wn_im[187] = $signed(16'sh5FE4);
  assign wn_im[188] = $signed(16'sh5ED7);
  assign wn_im[189] = $signed(16'sh5DC8);
  assign wn_im[190] = $signed(16'sh5CB4);
  assign wn_im[191] = $signed(16'sh5B9D);
  assign wn_im[192] = $signed(16'sh5A82);
  assign wn_im[193] = $signed(16'sh5964);
  assign wn_im[194] = $signed(16'sh5843);
  assign wn_im[195] = $signed(16'sh571E);
  assign wn_im[196] = $signed(16'sh55F6);
  assign wn_im[197] = $signed(16'sh54CA);
  assign wn_im[198] = $signed(16'sh539B);
  assign wn_im[199] = $signed(16'sh5269);
  assign wn_im[200] = $signed(16'sh5134);
  assign wn_im[201] = $signed(16'sh4FFB);
  assign wn_im[202] = $signed(16'sh4EC0);
  assign wn_im[203] = $signed(16'sh4D81);
  assign wn_im[204] = $signed(16'sh4C40);
  assign wn_im[205] = $signed(16'sh4AFB);
  assign wn_im[206] = $signed(16'sh49B4);
  assign wn_im[207] = $signed(16'sh486A);
  assign wn_im[208] = $signed(16'sh471D);
  assign wn_im[209] = $signed(16'sh45CD);
  assign wn_im[210] = $signed(16'sh447B);
  assign wn_im[211] = $signed(16'sh4326);
  assign wn_im[212] = $signed(16'sh41CE);
  assign wn_im[213] = $signed(16'sh4074);
  assign wn_im[214] = $signed(16'sh3F17);
  assign wn_im[215] = $signed(16'sh3DB8);
  assign wn_im[216] = $signed(16'sh3C57);
  assign wn_im[217] = $signed(16'sh3AF3);
  assign wn_im[218] = $signed(16'sh398D);
  assign wn_im[219] = $signed(16'sh3825);
  assign wn_im[220] = $signed(16'sh36BA);
  assign wn_im[221] = $signed(16'sh354E);
  assign wn_im[222] = $signed(16'sh33DF);
  assign wn_im[223] = $signed(16'sh326E);
  assign wn_im[224] = $signed(16'sh30FC);
  assign wn_im[225] = $signed(16'sh2F87);
  assign wn_im[226] = $signed(16'sh2E11);
  assign wn_im[227] = $signed(16'sh2C99);
  assign wn_im[228] = $signed(16'sh2B1F);
  assign wn_im[229] = $signed(16'sh29A4);
  assign wn_im[230] = $signed(16'sh2827);
  assign wn_im[231] = $signed(16'sh26A8);
  assign wn_im[232] = $signed(16'sh2528);
  assign wn_im[233] = $signed(16'sh23A7);
  assign wn_im[234] = $signed(16'sh2224);
  assign wn_im[235] = $signed(16'sh209F);
  assign wn_im[236] = $signed(16'sh1F1A);
  assign wn_im[237] = $signed(16'sh1D93);
  assign wn_im[238] = $signed(16'sh1C0C);
  assign wn_im[239] = $signed(16'sh1A83);
  assign wn_im[240] = $signed(16'sh18F9);
  assign wn_im[241] = $signed(16'sh176E);
  assign wn_im[242] = $signed(16'sh15E2);
  assign wn_im[243] = $signed(16'sh1455);
  assign wn_im[244] = $signed(16'sh12C8);
  assign wn_im[245] = $signed(16'sh113A);
  assign wn_im[246] = $signed(16'sh0FAB);
  assign wn_im[247] = $signed(16'sh0E1C);
  assign wn_im[248] = $signed(16'sh0C8C);
  assign wn_im[249] = $signed(16'sh0AFB);
  assign wn_im[250] = $signed(16'sh096B);
  assign wn_im[251] = $signed(16'sh07D9);
  assign wn_im[252] = $signed(16'sh0648);
  assign wn_im[253] = $signed(16'sh04B6);
  assign wn_im[254] = $signed(16'sh0324);
  assign wn_im[255] = $signed(16'sh0192);

  assign data0_re = wn_re[addr0];
  assign data0_im = wn_im[addr0];
  assign data1_re = wn_re[addr1];
  assign data1_im = wn_im[addr1];
  assign data2_re = wn_re[addr2];
  assign data2_im = wn_im[addr2];
  assign data3_re = wn_re[addr3];
  assign data3_im = wn_im[addr3];
  assign data4_re = wn_re[addr4];
  assign data4_im = wn_im[addr4];
  assign data5_re = wn_re[addr5];
  assign data5_im = wn_im[addr5];
  assign data6_re = wn_re[addr6];
  assign data6_im = wn_im[addr6];
  assign data7_re = wn_re[addr7];
  assign data7_im = wn_im[addr7];

endmodule  